// Code your testbench here
// or browse Examples
module mux_test();
  reg [7:0] bin1;
    reg [2:0]bctrl;
    wire bout;
        wire dum1,dum5;
  wire [3:0]dum2,dum6;
  wire [7:0] dum3,dum4;
    reg [31:0] data[0:2];
  initial $readmemh("lut_mux.mem",data);
    reg wclock;
    initial wclock=0;
    always #10 wclock=!wclock;
    FGPA ha_ha(.in1(bin1[7]),.in2(bin1[6]),.in3(bin1[5]),.in4(bin1[4]),.in5(bin1[3]),.in6(bin1[2]),.in7(bin1[1]),.in8(bin1[0]),.clock(wclock),.ctr1(bctrl[2]),.ctr2(bctrl[1]),.ctr3(bctrl[0]),.out(dum6),.out_carry(dum1),.sum_out(dum2),.q(dum3),.prev(dum4),.si(dum5),.out_mux(bout));
    initial
        begin
          ha_ha.l1.mem={data[1][0],data[2]};
          ha_ha.l2.mem={data[1][0],data[2]};
          ha_ha.l3.mem={data[1][0],data[2]};
          ha_ha.l4.mem={data[1][0],data[2]};
          ha_ha.l5.mem={data[1][0],data[2]};
          ha_ha.l6.mem={data[1][0],data[2]};
          ha_ha.l7.mem={data[1][0],data[2]};
          ha_ha.l8.mem={data[1][0],data[2]};
          ha_ha.l9.mem={data[1][0],data[2]};
          ha_ha.l10.mem={data[1][0],data[2]};
          ha_ha.l11.mem={data[1][0],data[2]};
          ha_ha.l12.mem={data[1][0],data[2]};
          ha_ha.l13.mem={data[1][0],data[2]};
          ha_ha.l14.mem={data[1][0],data[2]};
          ha_ha.l15.mem={data[1][0],data[2]};
          ha_ha.l16.mem={data[1][0],data[2]};
          ha_ha.l17.mem={data[1][0],data[2]};
            ha_ha.l18.mem={data[1][0],data[0]};
            ha_ha.l19.mem={data[1][0],data[0]};
            ha_ha.l20.mem={data[1][0],data[0]};
            ha_ha.l21.mem={data[1][0],data[0]};
            ha_ha.l22.mem={data[1][0],data[0]};
            ha_ha.l23.mem={data[1][0],data[0]};
            ha_ha.l24.mem={data[1][0],data[0]};
          ha_ha.l25.mem={data[1][0],data[2]};
          ha_ha.l26.mem={data[1][0],data[2]};
          ha_ha.l27.mem={data[1][0],data[2]};
          ha_ha.l28.mem={data[1][0],data[2]};
          ha_ha.l29.mem={data[1][0],data[2]};
          ha_ha.l30.mem={data[1][0],data[2]};
          ha_ha.l31.mem={data[1][0],data[2]};
          ha_ha.l32.mem={data[1][0],data[2]};
          ha_ha.l33.mem={data[1][0],data[2]};
          ha_ha.l34.mem={data[1][0],data[2]};
          ha_ha.l35.mem={data[1][0],data[2]};
          ha_ha.l36.mem={data[1][0],data[2]};
          ha_ha.l37.mem={data[1][0],data[2]};
          ha_ha.l38.mem={data[1][0],data[2]};
          ha_ha.l39.mem={data[1][0],data[2]};
          ha_ha.l40.mem={data[1][0],data[2]};
          ha_ha.l41.mem={data[1][0],data[2]};
          ha_ha.l42.mem={data[1][0],data[2]};
          ha_ha.l43.mem={data[1][0],data[2]};
          ha_ha.l44.mem={data[1][0],data[2]};
          ha_ha.l45.mem={data[1][0],data[2]};
          ha_ha.l46.mem={data[1][0],data[2]};
          ha_ha.l47.mem={data[1][0],data[2]};
          ha_ha.l48.mem={data[1][0],data[2]};
            bin1=8'b11010010;
            bctrl=3'b000;
            #10
            $display("%b",bout);

            ha_ha.l1.mem={data[1][0],data[2]};
          ha_ha.l2.mem={data[1][0],data[2]};
          ha_ha.l3.mem={data[1][0],data[2]};
          ha_ha.l4.mem={data[1][0],data[2]};
          ha_ha.l5.mem={data[1][0],data[2]};
          ha_ha.l6.mem={data[1][0],data[2]};
          ha_ha.l7.mem={data[1][0],data[2]};
          ha_ha.l8.mem={data[1][0],data[2]};
          ha_ha.l9.mem={data[1][0],data[2]};
          ha_ha.l10.mem={data[1][0],data[2]};
          ha_ha.l11.mem={data[1][0],data[2]};
          ha_ha.l12.mem={data[1][0],data[2]};
          ha_ha.l13.mem={data[1][0],data[2]};
          ha_ha.l14.mem={data[1][0],data[2]};
          ha_ha.l15.mem={data[1][0],data[2]};
          ha_ha.l16.mem={data[1][0],data[2]};
          ha_ha.l17.mem={data[1][0],data[2]};
            ha_ha.l18.mem={data[1][0],data[0]};
            ha_ha.l19.mem={data[1][0],data[0]};
            ha_ha.l20.mem={data[1][0],data[0]};
            ha_ha.l21.mem={data[1][0],data[0]};
            ha_ha.l22.mem={data[1][0],data[0]};
            ha_ha.l23.mem={data[1][0],data[0]};
            ha_ha.l24.mem={data[1][0],data[0]};
          ha_ha.l25.mem={data[1][0],data[2]};
          ha_ha.l26.mem={data[1][0],data[2]};
          ha_ha.l27.mem={data[1][0],data[2]};
          ha_ha.l28.mem={data[1][0],data[2]};
          ha_ha.l29.mem={data[1][0],data[2]};
          ha_ha.l30.mem={data[1][0],data[2]};
          ha_ha.l31.mem={data[1][0],data[2]};
          ha_ha.l32.mem={data[1][0],data[2]};
          ha_ha.l33.mem={data[1][0],data[2]};
          ha_ha.l34.mem={data[1][0],data[2]};
          ha_ha.l35.mem={data[1][0],data[2]};
          ha_ha.l36.mem={data[1][0],data[2]};
          ha_ha.l37.mem={data[1][0],data[2]};
          ha_ha.l38.mem={data[1][0],data[2]};
          ha_ha.l39.mem={data[1][0],data[2]};
          ha_ha.l40.mem={data[1][0],data[2]};
          ha_ha.l41.mem={data[1][0],data[2]};
          ha_ha.l42.mem={data[1][0],data[2]};
          ha_ha.l43.mem={data[1][0],data[2]};
          ha_ha.l44.mem={data[1][0],data[2]};
          ha_ha.l45.mem={data[1][0],data[2]};
          ha_ha.l46.mem={data[1][0],data[2]};
          ha_ha.l47.mem={data[1][0],data[2]};
          ha_ha.l48.mem={data[1][0],data[2]};
            bin1=8'b11010010;
            bctrl=3'b001;
            #10
            $display("%b",bout);

            ha_ha.l1.mem={data[1][0],data[2]};
          ha_ha.l2.mem={data[1][0],data[2]};
          ha_ha.l3.mem={data[1][0],data[2]};
          ha_ha.l4.mem={data[1][0],data[2]};
          ha_ha.l5.mem={data[1][0],data[2]};
          ha_ha.l6.mem={data[1][0],data[2]};
          ha_ha.l7.mem={data[1][0],data[2]};
          ha_ha.l8.mem={data[1][0],data[2]};
          ha_ha.l9.mem={data[1][0],data[2]};
          ha_ha.l10.mem={data[1][0],data[2]};
          ha_ha.l11.mem={data[1][0],data[2]};
          ha_ha.l12.mem={data[1][0],data[2]};
          ha_ha.l13.mem={data[1][0],data[2]};
          ha_ha.l14.mem={data[1][0],data[2]};
          ha_ha.l15.mem={data[1][0],data[2]};
          ha_ha.l16.mem={data[1][0],data[2]};
          ha_ha.l17.mem={data[1][0],data[2]};
            ha_ha.l18.mem={data[1][0],data[0]};
            ha_ha.l19.mem={data[1][0],data[0]};
            ha_ha.l20.mem={data[1][0],data[0]};
            ha_ha.l21.mem={data[1][0],data[0]};
            ha_ha.l22.mem={data[1][0],data[0]};
            ha_ha.l23.mem={data[1][0],data[0]};
            ha_ha.l24.mem={data[1][0],data[0]};
          ha_ha.l25.mem={data[1][0],data[2]};
          ha_ha.l26.mem={data[1][0],data[2]};
          ha_ha.l27.mem={data[1][0],data[2]};
          ha_ha.l28.mem={data[1][0],data[2]};
          ha_ha.l29.mem={data[1][0],data[2]};
          ha_ha.l30.mem={data[1][0],data[2]};
          ha_ha.l31.mem={data[1][0],data[2]};
          ha_ha.l32.mem={data[1][0],data[2]};
          ha_ha.l33.mem={data[1][0],data[2]};
          ha_ha.l34.mem={data[1][0],data[2]};
          ha_ha.l35.mem={data[1][0],data[2]};
          ha_ha.l36.mem={data[1][0],data[2]};
          ha_ha.l37.mem={data[1][0],data[2]};
          ha_ha.l38.mem={data[1][0],data[2]};
          ha_ha.l39.mem={data[1][0],data[2]};
          ha_ha.l40.mem={data[1][0],data[2]};
          ha_ha.l41.mem={data[1][0],data[2]};
          ha_ha.l42.mem={data[1][0],data[2]};
          ha_ha.l43.mem={data[1][0],data[2]};
          ha_ha.l44.mem={data[1][0],data[2]};
          ha_ha.l45.mem={data[1][0],data[2]};
          ha_ha.l46.mem={data[1][0],data[2]};
          ha_ha.l47.mem={data[1][0],data[2]};
          ha_ha.l48.mem={data[1][0],data[2]};
            bin1=8'b11010010;
            bctrl=3'b010;
            #10
            $display("%b",bout);

           ha_ha.l1.mem={data[1][0],data[2]};
          ha_ha.l2.mem={data[1][0],data[2]};
          ha_ha.l3.mem={data[1][0],data[2]};
          ha_ha.l4.mem={data[1][0],data[2]};
          ha_ha.l5.mem={data[1][0],data[2]};
          ha_ha.l6.mem={data[1][0],data[2]};
          ha_ha.l7.mem={data[1][0],data[2]};
          ha_ha.l8.mem={data[1][0],data[2]};
          ha_ha.l9.mem={data[1][0],data[2]};
          ha_ha.l10.mem={data[1][0],data[2]};
          ha_ha.l11.mem={data[1][0],data[2]};
          ha_ha.l12.mem={data[1][0],data[2]};
          ha_ha.l13.mem={data[1][0],data[2]};
          ha_ha.l14.mem={data[1][0],data[2]};
          ha_ha.l15.mem={data[1][0],data[2]};
          ha_ha.l16.mem={data[1][0],data[2]};
          ha_ha.l17.mem={data[1][0],data[2]};
            ha_ha.l18.mem={data[1][0],data[0]};
            ha_ha.l19.mem={data[1][0],data[0]};
            ha_ha.l20.mem={data[1][0],data[0]};
            ha_ha.l21.mem={data[1][0],data[0]};
            ha_ha.l22.mem={data[1][0],data[0]};
            ha_ha.l23.mem={data[1][0],data[0]};
            ha_ha.l24.mem={data[1][0],data[0]};
          ha_ha.l25.mem={data[1][0],data[2]};
          ha_ha.l26.mem={data[1][0],data[2]};
          ha_ha.l27.mem={data[1][0],data[2]};
          ha_ha.l28.mem={data[1][0],data[2]};
          ha_ha.l29.mem={data[1][0],data[2]};
          ha_ha.l30.mem={data[1][0],data[2]};
          ha_ha.l31.mem={data[1][0],data[2]};
          ha_ha.l32.mem={data[1][0],data[2]};
          ha_ha.l33.mem={data[1][0],data[2]};
          ha_ha.l34.mem={data[1][0],data[2]};
          ha_ha.l35.mem={data[1][0],data[2]};
          ha_ha.l36.mem={data[1][0],data[2]};
          ha_ha.l37.mem={data[1][0],data[2]};
          ha_ha.l38.mem={data[1][0],data[2]};
          ha_ha.l39.mem={data[1][0],data[2]};
          ha_ha.l40.mem={data[1][0],data[2]};
          ha_ha.l41.mem={data[1][0],data[2]};
          ha_ha.l42.mem={data[1][0],data[2]};
          ha_ha.l43.mem={data[1][0],data[2]};
          ha_ha.l44.mem={data[1][0],data[2]};
          ha_ha.l45.mem={data[1][0],data[2]};
          ha_ha.l46.mem={data[1][0],data[2]};
          ha_ha.l47.mem={data[1][0],data[2]};
          ha_ha.l48.mem={data[1][0],data[2]};
            bin1=8'b11010010;
            bctrl=3'b011;
            #10
            $display("%b",bout);

            ha_ha.l1.mem={data[1][0],data[2]};
          ha_ha.l2.mem={data[1][0],data[2]};
          ha_ha.l3.mem={data[1][0],data[2]};
          ha_ha.l4.mem={data[1][0],data[2]};
          ha_ha.l5.mem={data[1][0],data[2]};
          ha_ha.l6.mem={data[1][0],data[2]};
          ha_ha.l7.mem={data[1][0],data[2]};
          ha_ha.l8.mem={data[1][0],data[2]};
          ha_ha.l9.mem={data[1][0],data[2]};
          ha_ha.l10.mem={data[1][0],data[2]};
          ha_ha.l11.mem={data[1][0],data[2]};
          ha_ha.l12.mem={data[1][0],data[2]};
          ha_ha.l13.mem={data[1][0],data[2]};
          ha_ha.l14.mem={data[1][0],data[2]};
          ha_ha.l15.mem={data[1][0],data[2]};
          ha_ha.l16.mem={data[1][0],data[2]};
          ha_ha.l17.mem={data[1][0],data[2]};
            ha_ha.l18.mem={data[1][0],data[0]};
            ha_ha.l19.mem={data[1][0],data[0]};
            ha_ha.l20.mem={data[1][0],data[0]};
            ha_ha.l21.mem={data[1][0],data[0]};
            ha_ha.l22.mem={data[1][0],data[0]};
            ha_ha.l23.mem={data[1][0],data[0]};
            ha_ha.l24.mem={data[1][0],data[0]};
          ha_ha.l25.mem={data[1][0],data[2]};
          ha_ha.l26.mem={data[1][0],data[2]};
          ha_ha.l27.mem={data[1][0],data[2]};
          ha_ha.l28.mem={data[1][0],data[2]};
          ha_ha.l29.mem={data[1][0],data[2]};
          ha_ha.l30.mem={data[1][0],data[2]};
          ha_ha.l31.mem={data[1][0],data[2]};
          ha_ha.l32.mem={data[1][0],data[2]};
          ha_ha.l33.mem={data[1][0],data[2]};
          ha_ha.l34.mem={data[1][0],data[2]};
          ha_ha.l35.mem={data[1][0],data[2]};
          ha_ha.l36.mem={data[1][0],data[2]};
          ha_ha.l37.mem={data[1][0],data[2]};
          ha_ha.l38.mem={data[1][0],data[2]};
          ha_ha.l39.mem={data[1][0],data[2]};
          ha_ha.l40.mem={data[1][0],data[2]};
          ha_ha.l41.mem={data[1][0],data[2]};
          ha_ha.l42.mem={data[1][0],data[2]};
          ha_ha.l43.mem={data[1][0],data[2]};
          ha_ha.l44.mem={data[1][0],data[2]};
          ha_ha.l45.mem={data[1][0],data[2]};
          ha_ha.l46.mem={data[1][0],data[2]};
          ha_ha.l47.mem={data[1][0],data[2]};
          ha_ha.l48.mem={data[1][0],data[2]};
            bin1=8'b11010010;
            bctrl=3'b100;
            #10
            $display("%b",bout);

            ha_ha.l1.mem={data[1][0],data[2]};
          ha_ha.l2.mem={data[1][0],data[2]};
          ha_ha.l3.mem={data[1][0],data[2]};
          ha_ha.l4.mem={data[1][0],data[2]};
          ha_ha.l5.mem={data[1][0],data[2]};
          ha_ha.l6.mem={data[1][0],data[2]};
          ha_ha.l7.mem={data[1][0],data[2]};
          ha_ha.l8.mem={data[1][0],data[2]};
          ha_ha.l9.mem={data[1][0],data[2]};
          ha_ha.l10.mem={data[1][0],data[2]};
          ha_ha.l11.mem={data[1][0],data[2]};
          ha_ha.l12.mem={data[1][0],data[2]};
          ha_ha.l13.mem={data[1][0],data[2]};
          ha_ha.l14.mem={data[1][0],data[2]};
          ha_ha.l15.mem={data[1][0],data[2]};
          ha_ha.l16.mem={data[1][0],data[2]};
          ha_ha.l17.mem={data[1][0],data[2]};
            ha_ha.l18.mem={data[1][0],data[0]};
            ha_ha.l19.mem={data[1][0],data[0]};
            ha_ha.l20.mem={data[1][0],data[0]};
            ha_ha.l21.mem={data[1][0],data[0]};
            ha_ha.l22.mem={data[1][0],data[0]};
            ha_ha.l23.mem={data[1][0],data[0]};
            ha_ha.l24.mem={data[1][0],data[0]};
          ha_ha.l25.mem={data[1][0],data[2]};
          ha_ha.l26.mem={data[1][0],data[2]};
          ha_ha.l27.mem={data[1][0],data[2]};
          ha_ha.l28.mem={data[1][0],data[2]};
          ha_ha.l29.mem={data[1][0],data[2]};
          ha_ha.l30.mem={data[1][0],data[2]};
          ha_ha.l31.mem={data[1][0],data[2]};
          ha_ha.l32.mem={data[1][0],data[2]};
          ha_ha.l33.mem={data[1][0],data[2]};
          ha_ha.l34.mem={data[1][0],data[2]};
          ha_ha.l35.mem={data[1][0],data[2]};
          ha_ha.l36.mem={data[1][0],data[2]};
          ha_ha.l37.mem={data[1][0],data[2]};
          ha_ha.l38.mem={data[1][0],data[2]};
          ha_ha.l39.mem={data[1][0],data[2]};
          ha_ha.l40.mem={data[1][0],data[2]};
          ha_ha.l41.mem={data[1][0],data[2]};
          ha_ha.l42.mem={data[1][0],data[2]};
          ha_ha.l43.mem={data[1][0],data[2]};
          ha_ha.l44.mem={data[1][0],data[2]};
          ha_ha.l45.mem={data[1][0],data[2]};
          ha_ha.l46.mem={data[1][0],data[2]};
          ha_ha.l47.mem={data[1][0],data[2]};
          ha_ha.l48.mem={data[1][0],data[2]};
            bin1=8'b11010010;
            bctrl=3'b101;
            #10
            $display("%b",bout);

            ha_ha.l1.mem={data[1][0],data[2]};
          ha_ha.l2.mem={data[1][0],data[2]};
          ha_ha.l3.mem={data[1][0],data[2]};
          ha_ha.l4.mem={data[1][0],data[2]};
          ha_ha.l5.mem={data[1][0],data[2]};
          ha_ha.l6.mem={data[1][0],data[2]};
          ha_ha.l7.mem={data[1][0],data[2]};
          ha_ha.l8.mem={data[1][0],data[2]};
          ha_ha.l9.mem={data[1][0],data[2]};
          ha_ha.l10.mem={data[1][0],data[2]};
          ha_ha.l11.mem={data[1][0],data[2]};
          ha_ha.l12.mem={data[1][0],data[2]};
          ha_ha.l13.mem={data[1][0],data[2]};
          ha_ha.l14.mem={data[1][0],data[2]};
          ha_ha.l15.mem={data[1][0],data[2]};
          ha_ha.l16.mem={data[1][0],data[2]};
          ha_ha.l17.mem={data[1][0],data[2]};
            ha_ha.l18.mem={data[1][0],data[0]};
            ha_ha.l19.mem={data[1][0],data[0]};
            ha_ha.l20.mem={data[1][0],data[0]};
            ha_ha.l21.mem={data[1][0],data[0]};
            ha_ha.l22.mem={data[1][0],data[0]};
            ha_ha.l23.mem={data[1][0],data[0]};
            ha_ha.l24.mem={data[1][0],data[0]};
          ha_ha.l25.mem={data[1][0],data[2]};
          ha_ha.l26.mem={data[1][0],data[2]};
          ha_ha.l27.mem={data[1][0],data[2]};
          ha_ha.l28.mem={data[1][0],data[2]};
          ha_ha.l29.mem={data[1][0],data[2]};
          ha_ha.l30.mem={data[1][0],data[2]};
          ha_ha.l31.mem={data[1][0],data[2]};
          ha_ha.l32.mem={data[1][0],data[2]};
          ha_ha.l33.mem={data[1][0],data[2]};
          ha_ha.l34.mem={data[1][0],data[2]};
          ha_ha.l35.mem={data[1][0],data[2]};
          ha_ha.l36.mem={data[1][0],data[2]};
          ha_ha.l37.mem={data[1][0],data[2]};
          ha_ha.l38.mem={data[1][0],data[2]};
          ha_ha.l39.mem={data[1][0],data[2]};
          ha_ha.l40.mem={data[1][0],data[2]};
          ha_ha.l41.mem={data[1][0],data[2]};
          ha_ha.l42.mem={data[1][0],data[2]};
          ha_ha.l43.mem={data[1][0],data[2]};
          ha_ha.l44.mem={data[1][0],data[2]};
          ha_ha.l45.mem={data[1][0],data[2]};
          ha_ha.l46.mem={data[1][0],data[2]};
          ha_ha.l47.mem={data[1][0],data[2]};
          ha_ha.l48.mem={data[1][0],data[2]};
            bin1=8'b11010010;
            bctrl=3'b110;
            #10
            $display("%b",bout);

            ha_ha.l1.mem={data[1][0],data[2]};
          ha_ha.l2.mem={data[1][0],data[2]};
          ha_ha.l3.mem={data[1][0],data[2]};
          ha_ha.l4.mem={data[1][0],data[2]};
          ha_ha.l5.mem={data[1][0],data[2]};
          ha_ha.l6.mem={data[1][0],data[2]};
          ha_ha.l7.mem={data[1][0],data[2]};
          ha_ha.l8.mem={data[1][0],data[2]};
          ha_ha.l9.mem={data[1][0],data[2]};
          ha_ha.l10.mem={data[1][0],data[2]};
          ha_ha.l11.mem={data[1][0],data[2]};
          ha_ha.l12.mem={data[1][0],data[2]};
          ha_ha.l13.mem={data[1][0],data[2]};
          ha_ha.l14.mem={data[1][0],data[2]};
          ha_ha.l15.mem={data[1][0],data[2]};
          ha_ha.l16.mem={data[1][0],data[2]};
          ha_ha.l17.mem={data[1][0],data[2]};
            ha_ha.l18.mem={data[1][0],data[0]};
            ha_ha.l19.mem={data[1][0],data[0]};
            ha_ha.l20.mem={data[1][0],data[0]};
            ha_ha.l21.mem={data[1][0],data[0]};
            ha_ha.l22.mem={data[1][0],data[0]};
            ha_ha.l23.mem={data[1][0],data[0]};
            ha_ha.l24.mem={data[1][0],data[0]};
          ha_ha.l25.mem={data[1][0],data[2]};
          ha_ha.l26.mem={data[1][0],data[2]};
          ha_ha.l27.mem={data[1][0],data[2]};
          ha_ha.l28.mem={data[1][0],data[2]};
          ha_ha.l29.mem={data[1][0],data[2]};
          ha_ha.l30.mem={data[1][0],data[2]};
          ha_ha.l31.mem={data[1][0],data[2]};
          ha_ha.l32.mem={data[1][0],data[2]};
          ha_ha.l33.mem={data[1][0],data[2]};
          ha_ha.l34.mem={data[1][0],data[2]};
          ha_ha.l35.mem={data[1][0],data[2]};
          ha_ha.l36.mem={data[1][0],data[2]};
          ha_ha.l37.mem={data[1][0],data[2]};
          ha_ha.l38.mem={data[1][0],data[2]};
          ha_ha.l39.mem={data[1][0],data[2]};
          ha_ha.l40.mem={data[1][0],data[2]};
          ha_ha.l41.mem={data[1][0],data[2]};
          ha_ha.l42.mem={data[1][0],data[2]};
          ha_ha.l43.mem={data[1][0],data[2]};
          ha_ha.l44.mem={data[1][0],data[2]};
          ha_ha.l45.mem={data[1][0],data[2]};
          ha_ha.l46.mem={data[1][0],data[2]};
          ha_ha.l47.mem={data[1][0],data[2]};
          ha_ha.l48.mem={data[1][0],data[2]};
            bin1=8'b11010010;
            bctrl=3'b111;
            #10
            $display("%b",bout);

            $finish;
        end
    initial
        begin
          $dumpfile("ha_mux.vcd");
            $dumpvars;
        end
endmodule


module switch_test();
    reg [7:0] bin1;
    reg [2:0]bctrl;
    wire bout;
        wire dum1;
  reg rsi;
  wire [3:0]dum2,dum6;
  wire [7:0] rq;
  reg [7:0]rprev;
  initial rprev=8'b00000000;
  always #15 rprev=rq;
    reg [31:0] data[0:2];
  initial $readmemh("lut_register.mem",data);
    reg wclock;
    initial wclock=0;
    always #10 wclock=!wclock;
    FGPA ha_ha(.in1(bin1[7]),.in2(bin1[6]),.in3(bin1[5]),.in4(bin1[4]),.in5(bin1[3]),.in6(bin1[2]),.in7(bin1[1]),.in8(bin1[0]),.clock(wclock),.ctr1(bctrl[2]),.ctr2(bctrl[1]),.ctr3(bctrl[0]),.out(dum6),.out_carry(dum1),.sum_out(dum2),.q(rq),.prev(rprev),.si(rsi),.out_mux(bout));
    initial
        begin
            ha_ha.l1.mem={data[1][0],data[2]};
          ha_ha.l2.mem={data[1][0],data[2]};
          ha_ha.l3.mem={data[1][0],data[2]};
          ha_ha.l4.mem={data[1][0],data[2]};
          ha_ha.l5.mem={data[1][0],data[2]};
          ha_ha.l6.mem={data[1][0],data[2]};
          ha_ha.l7.mem={data[1][0],data[2]};
          ha_ha.l8.mem={data[1][0],data[2]};
          ha_ha.l9.mem={data[1][0],data[2]};
          ha_ha.l10.mem={data[1][0],data[2]};
          ha_ha.l11.mem={data[1][0],data[2]};
          ha_ha.l12.mem={data[1][0],data[2]};
          ha_ha.l13.mem={data[1][0],data[2]};
          ha_ha.l14.mem={data[1][0],data[2]};
          ha_ha.l15.mem={data[1][0],data[2]};
          ha_ha.l16.mem={data[1][0],data[2]};
          ha_ha.l17.mem={data[1][0],data[2]};
          ha_ha.l18.mem={data[1][0],data[2]};
          ha_ha.l19.mem={data[1][0],data[2]};
          ha_ha.l20.mem={data[1][0],data[2]};
          ha_ha.l21.mem={data[1][0],data[2]};
          ha_ha.l22.mem={data[1][0],data[2]};
          ha_ha.l23.mem={data[1][0],data[2]};
          ha_ha.l24.mem={data[1][0],data[2]};
          ha_ha.l25.mem={data[1][0],data[0]};
          ha_ha.l26.mem={data[1][0],data[0]};
          ha_ha.l27.mem={data[1][0],data[0]};
          ha_ha.l28.mem={data[1][0],data[0]};
          ha_ha.l29.mem={data[1][0],data[0]};
          ha_ha.l30.mem={data[1][0],data[0]};
          ha_ha.l31.mem={data[1][0],data[0]};
          ha_ha.l32.mem={data[1][0],data[0]};
          ha_ha.l33.mem={data[1][0],data[0]};
          ha_ha.l34.mem={data[1][0],data[0]};
          ha_ha.l35.mem={data[1][0],data[0]};
          ha_ha.l36.mem={data[1][0],data[0]};
          ha_ha.l37.mem={data[1][0],data[0]};
          ha_ha.l38.mem={data[1][0],data[0]};
          ha_ha.l39.mem={data[1][0],data[0]};
          ha_ha.l40.mem={data[1][0],data[0]};
          ha_ha.l41.mem={data[1][0],data[0]};
          ha_ha.l42.mem={data[1][0],data[0]};
          ha_ha.l43.mem={data[1][0],data[0]};
          ha_ha.l44.mem={data[1][0],data[0]};
          ha_ha.l45.mem={data[1][0],data[0]};
          ha_ha.l46.mem={data[1][0],data[0]};
          ha_ha.l47.mem={data[1][0],data[0]};
          ha_ha.l48.mem={data[1][0],data[0]};
            bin1=8'b10110010;
            rsi=1'b1;
            bctrl=3'b001;
          #15
          $display("%b",rq);

          ha_ha.l1.mem={data[1][0],data[2]};
          ha_ha.l2.mem={data[1][0],data[2]};
          ha_ha.l3.mem={data[1][0],data[2]};
          ha_ha.l4.mem={data[1][0],data[2]};
          ha_ha.l5.mem={data[1][0],data[2]};
          ha_ha.l6.mem={data[1][0],data[2]};
          ha_ha.l7.mem={data[1][0],data[2]};
          ha_ha.l8.mem={data[1][0],data[2]};
          ha_ha.l9.mem={data[1][0],data[2]};
          ha_ha.l10.mem={data[1][0],data[2]};
          ha_ha.l11.mem={data[1][0],data[2]};
          ha_ha.l12.mem={data[1][0],data[2]};
          ha_ha.l13.mem={data[1][0],data[2]};
          ha_ha.l14.mem={data[1][0],data[2]};
          ha_ha.l15.mem={data[1][0],data[2]};
          ha_ha.l16.mem={data[1][0],data[2]};
          ha_ha.l17.mem={data[1][0],data[2]};
          ha_ha.l18.mem={data[1][0],data[2]};
          ha_ha.l19.mem={data[1][0],data[2]};
          ha_ha.l20.mem={data[1][0],data[2]};
          ha_ha.l21.mem={data[1][0],data[2]};
          ha_ha.l22.mem={data[1][0],data[2]};
          ha_ha.l23.mem={data[1][0],data[2]};
          ha_ha.l24.mem={data[1][0],data[2]};
          ha_ha.l25.mem={data[1][0],data[0]};
          ha_ha.l26.mem={data[1][0],data[0]};
          ha_ha.l27.mem={data[1][0],data[0]};
          ha_ha.l28.mem={data[1][0],data[0]};
          ha_ha.l29.mem={data[1][0],data[0]};
          ha_ha.l30.mem={data[1][0],data[0]};
          ha_ha.l31.mem={data[1][0],data[0]};
          ha_ha.l32.mem={data[1][0],data[0]};
          ha_ha.l33.mem={data[1][0],data[0]};
          ha_ha.l34.mem={data[1][0],data[0]};
          ha_ha.l35.mem={data[1][0],data[0]};
          ha_ha.l36.mem={data[1][0],data[0]};
          ha_ha.l37.mem={data[1][0],data[0]};
          ha_ha.l38.mem={data[1][0],data[0]};
          ha_ha.l39.mem={data[1][0],data[0]};
          ha_ha.l40.mem={data[1][0],data[0]};
          ha_ha.l41.mem={data[1][0],data[0]};
          ha_ha.l42.mem={data[1][0],data[0]};
          ha_ha.l43.mem={data[1][0],data[0]};
          ha_ha.l44.mem={data[1][0],data[0]};
          ha_ha.l45.mem={data[1][0],data[0]};
          ha_ha.l46.mem={data[1][0],data[0]};
          ha_ha.l47.mem={data[1][0],data[0]};
          ha_ha.l48.mem={data[1][0],data[0]};
            bin1=8'b10110010;
            rsi=1'b1;
            bctrl=3'b010;
          #15
          $display("%b",rq);
            $finish;
        end
endmodule



module bcd_test();
  reg [7:0] bin1;
    reg [2:0]bctrl;
    wire bout;
        wire dum1;
  wire rsi;
  wire [3:0]dum2,bcd_out;
  wire [7:0] rq;
  wire [7:0]rprev;
  reg [31:0] data[0:3
                 ];
  initial $readmemh("lut_bcd.mem",data);
    reg wclock;
    initial wclock=0;
    always #10 wclock=!wclock;
    FGPA ha_ha(.in1(bin1[7]),.in2(bin1[6]),.in3(bin1[5]),.in4(bin1[4]),.in5(bin1[3]),.in6(bin1[2]),.in7(bin1[1]),.in8(bin1[0]),.clock(wclock),.ctr1(bctrl[2]),.ctr2(bctrl[1]),.ctr3(bctrl[0]),.out(bcd_out),.out_carry(dum1),.sum_out(dum2),.q(rq),.prev(rprev),.si(rsi),.out_mux(bout));
  initial
        begin
            ha_ha.l1.mem={data[1][0],data[2]};
          ha_ha.l2.mem={data[1][0],data[2]};
          ha_ha.l3.mem={data[1][0],data[2]};
          ha_ha.l4.mem={data[1][0],data[2]};
          ha_ha.l5.mem={data[1][0],data[2]};
          ha_ha.l6.mem={data[1][0],data[2]};
          ha_ha.l7.mem={data[1][0],data[2]};
          ha_ha.l8.mem={data[1][0],data[2]};
          ha_ha.l9.mem={data[1][0],data[3]};
          ha_ha.l10.mem={data[1][0],data[2]};
          ha_ha.l11.mem={data[1][0],data[2]};
          ha_ha.l12.mem={data[1][0],data[2]};
          ha_ha.l13.mem={data[1][0],data[2]};
          ha_ha.l14.mem={data[1][0],data[2]};
          ha_ha.l15.mem={data[1][0],data[2]};
          ha_ha.l16.mem={data[1][0],data[2]};
          ha_ha.l17.mem={data[1][0],data[2]};
          ha_ha.l18.mem={data[1][0],data[0]};
          ha_ha.l19.mem={data[1][0],data[0]};
          ha_ha.l20.mem={data[1][0],data[0]};
          ha_ha.l21.mem={data[1][0],data[0]};
          ha_ha.l22.mem={data[1][0],data[0]};
          ha_ha.l23.mem={data[1][0],data[0]};
          ha_ha.l24.mem={data[1][0],data[0]};
          ha_ha.l25.mem={data[1][0],data[0]};
          ha_ha.l26.mem={data[1][0],data[0]};
          ha_ha.l27.mem={data[1][0],data[0]};
          ha_ha.l28.mem={data[1][0],data[0]};
          ha_ha.l29.mem={data[1][0],data[0]};
          ha_ha.l30.mem={data[1][0],data[0]};
          ha_ha.l31.mem={data[1][0],data[0]};
          ha_ha.l32.mem={data[1][0],data[0]};
          ha_ha.l33.mem={data[1][0],data[0]};
          ha_ha.l34.mem={data[1][0],data[0]};
          ha_ha.l35.mem={data[1][0],data[0]};
          ha_ha.l36.mem={data[1][0],data[0]};
          ha_ha.l37.mem={data[1][0],data[0]};
          ha_ha.l38.mem={data[1][0],data[0]};
          ha_ha.l39.mem={data[1][0],data[0]};
          ha_ha.l40.mem={data[1][0],data[0]};
          ha_ha.l41.mem={data[1][0],data[0]};
          ha_ha.l42.mem={data[1][0],data[0]};
          ha_ha.l43.mem={data[1][0],data[0]};
          ha_ha.l44.mem={data[1][0],data[0]};
          ha_ha.l45.mem={data[1][0],data[0]};
          ha_ha.l46.mem={data[1][0],data[0]};
          ha_ha.l47.mem={data[1][0],data[0]};
          ha_ha.l48.mem={data[1][0],data[0]};
            bin1=8'b10110010;
          bctrl[2]=1'b1;
          #10
          $display("%b %b",bcd_out,dum1);

          ha_ha.l1.mem={data[1][0],data[2]};
          ha_ha.l2.mem={data[1][0],data[2]};
          ha_ha.l3.mem={data[1][0],data[2]};
          ha_ha.l4.mem={data[1][0],data[2]};
          ha_ha.l5.mem={data[1][0],data[2]};
          ha_ha.l6.mem={data[1][0],data[2]};
          ha_ha.l7.mem={data[1][0],data[2]};
          ha_ha.l8.mem={data[1][0],data[2]};
          ha_ha.l9.mem={data[1][0],data[3]};
          ha_ha.l10.mem={data[1][0],data[2]};
          ha_ha.l11.mem={data[1][0],data[2]};
          ha_ha.l12.mem={data[1][0],data[2]};
          ha_ha.l13.mem={data[1][0],data[2]};
          ha_ha.l14.mem={data[1][0],data[2]};
          ha_ha.l15.mem={data[1][0],data[2]};
          ha_ha.l16.mem={data[1][0],data[2]};
          ha_ha.l17.mem={data[1][0],data[2]};
          ha_ha.l18.mem={data[1][0],data[0]};
          ha_ha.l19.mem={data[1][0],data[0]};
          ha_ha.l20.mem={data[1][0],data[0]};
          ha_ha.l21.mem={data[1][0],data[0]};
          ha_ha.l22.mem={data[1][0],data[0]};
          ha_ha.l23.mem={data[1][0],data[0]};
          ha_ha.l24.mem={data[1][0],data[0]};
          ha_ha.l25.mem={data[1][0],data[0]};
          ha_ha.l26.mem={data[1][0],data[0]};
          ha_ha.l27.mem={data[1][0],data[0]};
          ha_ha.l28.mem={data[1][0],data[0]};
          ha_ha.l29.mem={data[1][0],data[0]};
          ha_ha.l30.mem={data[1][0],data[0]};
          ha_ha.l31.mem={data[1][0],data[0]};
          ha_ha.l32.mem={data[1][0],data[0]};
          ha_ha.l33.mem={data[1][0],data[0]};
          ha_ha.l34.mem={data[1][0],data[0]};
          ha_ha.l35.mem={data[1][0],data[0]};
          ha_ha.l36.mem={data[1][0],data[0]};
          ha_ha.l37.mem={data[1][0],data[0]};
          ha_ha.l38.mem={data[1][0],data[0]};
          ha_ha.l39.mem={data[1][0],data[0]};
          ha_ha.l40.mem={data[1][0],data[0]};
          ha_ha.l41.mem={data[1][0],data[0]};
          ha_ha.l42.mem={data[1][0],data[0]};
          ha_ha.l43.mem={data[1][0],data[0]};
          ha_ha.l44.mem={data[1][0],data[0]};
          ha_ha.l45.mem={data[1][0],data[0]};
          ha_ha.l46.mem={data[1][0],data[0]};
          ha_ha.l47.mem={data[1][0],data[0]};
          ha_ha.l48.mem={data[1][0],data[0]};
            bin1=8'b11111010;
          bctrl[2]=1'b1;
          #10
          $display("%b %b",bcd_out,dum1);

        end
endmodule
